module current_monitor();

endmodule

