module sensor_position();

endmodule

