module control_pid();


endmodule

