module sensor_reader();

endmodule

